module hello_world();
  display("hello world");
endmodule
